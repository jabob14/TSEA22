library ieee;
  use ieee.std_logic_1164.all;

entity enpulsare is
  port (
    clk : in  std_logic;
    x   : in  std_logic;
    u   : out std_logic
  );
end entity;

architecture behav of enpulsare is
begin

end architecture;

